`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// 
//////////////////////////////////////////////////////////////////////////////////


module formula_test(
    output wire [33:0] out
    );
    
   parameter out1 = (1-2*3.14159265/10000000*10000)*67108864;
   assign out = out1;
    
endmodule
