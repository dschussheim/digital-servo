`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    14:24:29 06/01/2017 
// Design Name: 
// Module Name:    DAC_const_test 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//	Module to test if we can see constant values out of DAC.
//
//////////////////////////////////////////////////////////////////////////////////
module DAC_const_test(
    input [15:0] DAC1_in,
    input [15:0] DAC2_in,
    input clk_in,
    input [15:0] D_out_p,
    input [15:0] D_out_n
    );


endmodule
